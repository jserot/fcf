library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library fcf;
use fcf.utils.all;
use fcf.values.all;

package types is
  type r_arr32 is array(0 to 31) of real;
end package;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library fcf;
use fcf.utils.all;
use fcf.values.all;

use work.types.all;
package consts is
  constant x0: r_arr32;
  constant arctan: r_arr32;
end package;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library fcf;
use fcf.utils.all;
use fcf.values.all;

package body consts is
  constant x0: r_arr32 := (0.707106781187,0.632455532034,0.613571991078,0.608833912518,0.607648256256,0.607351770141,0.607277644094,0.607259112299,0.607254479333,0.60725332109,0.607253031529,0.607252959139,0.607252941041,0.607252936517,0.607252935386,0.607252935103,0.607252935032,0.607252935015,0.60725293501,0.607252935009,0.607252935009,0.607252935009,0.607252935009,0.607252935009,0.607252935009,0.607252935009,0.607252935009,0.607252935009,0.607252935009,0.607252935009,0.607252935009,0.607252935009);
  constant arctan: r_arr32 := (45.0,26.5650511771,14.0362434679,7.1250163489,3.576334375,1.78991060825,0.895173710211,0.447614170861,0.223810500369,0.111905677066,0.0559528918938,0.027976452617,0.0139882271423,0.00699411367535,0.0034970568507,0.00174852842698,0.000874264213694,0.000437132106872,0.000218566053439,0.00010928302672,5.46415133601e-05,2.732075668e-05,1.366037834e-05,6.83018917e-06,3.415094585e-06,1.7075472925e-06,8.537736463e-07,4.268868231e-07,2.134434116e-07,1.067217058e-07,5.33608529e-08,2.66804264e-08);
end package body;
